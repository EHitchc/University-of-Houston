** Profile: "SCHEMATIC1-Test"  [ C:\Users\Ethan\Documents\ECE 3456\Lab 5\Step A\cmos transmission gate-pspicefiles\schematic1\test.sim ] 

** Creating circuit file "Test.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../cmos transmission gate-PSpiceFiles/2input nand enhancement load.lib" 
.LIB "../../../cmos transmission gate-PSpiceFiles/2INPUT NOR ENHANCEMENT LOAD.lib" 
* From [PSPICE NETLIST] section of C:\Users\Ethan\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_A 0 5 1 
+ LIN V_Vin 0 5 1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
