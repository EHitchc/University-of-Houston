** Profile: "SCHEMATIC1-Test"  [ c:\users\ethan\documents\ece 3456\lab 4\step b - nand\2input nand cmos-PSpiceFiles\SCHEMATIC1\Test.sim ] 

** Creating circuit file "Test.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../2input nand cmos-PSpiceFiles/2INPUT NOR CMOS.lib" 
.LIB "../../../2input nand cmos-PSpiceFiles/2INPUT NOR ENHANCEMENT LOAD.lib" 
* From [PSPICE NETLIST] section of C:\Users\Ethan\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
